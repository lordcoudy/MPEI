* \\vmware-host\Shared Folders\�����������\LR_03 DO\LR3 1PP_1C.sch

* Schematics Version 9.2
* Mon Mar 22 15:03:57 2021



** Analysis setup **
.tran 10ns 2.4m 0.8m 0.8u
.four 1250 3 v([2])


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "LR3 1PP_1C.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
