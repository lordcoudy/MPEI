* \\vmware-host\Shared Folders\�����������\LR_03 DO\LR3 BAX_stab.sch

* Schematics Version 9.2
* Mon Mar 22 16:32:54 2021



** Analysis setup **
.DC LIN I_I1 -20m 20m 50u 
.LIB "C:\Diodes.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "LR3 BAX_stab.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
