* \\vmware-host\Shared Folders\�����������\LR_03 DO\LR3 2SO.sch

* Schematics Version 9.2
* Mon Mar 22 15:50:40 2021



** Analysis setup **
.tran 10ns 2m 0 3u
.LIB "C:\Diodes.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "LR3 2SO.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
