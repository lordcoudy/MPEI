* \\vmware-host\Shared Folders\�����������\LR_04 DO\BAX_OE.sch

* Schematics Version 9.2
* Tue Apr 13 14:54:33 2021



** Analysis setup **
.DC LIN V_V1 0 10 50m 
+ LIN I_I1 20u 300u 20u 
.LIB "C:\KP_2021\bipolar.lib"
.LIB "C:\KP_2021\RUS_Q.LIB"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "BAX_OE.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
