* C:\KP_2021\BAX_OE.sch

* Schematics Version 9.2
* Mon May 03 13:17:26 2021



** Analysis setup **
.DC LIN V_V1 0 40 15m 
+ LIN I_I1 50u 500u 50u 
.LIB "C:\KP_2021\bipolar.lib"
.LIB "C:\KP_2021\RUS_Q.LIB"
.LIB "C:\Diodes.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "BAX_OE.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
