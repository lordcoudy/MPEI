* C:\KP_2021\BAX_OE_V_yurach.sch

* Schematics Version 9.2
* Tue Apr 27 19:17:41 2021



** Analysis setup **
.DC LIN I_I1 0 500u 10n 
.LIB "C:\KP_2021\bipolar.lib"
.LIB "C:\KP_2021\RUS_Q.LIB"
.LIB "C:\Diodes.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "BAX_OE_V_yurach.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
