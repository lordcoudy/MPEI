* C:\KP_2021\RT.sch

* Schematics Version 9.2
* Sat May 08 14:32:37 2021



** Analysis setup **
.OP 
.LIB "C:\KP_2021\bipolar.lib"
.LIB "C:\KP_2021\Diodes.lib"
.LIB "C:\KP_2021\RUS_Q.LIB"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "RT.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
